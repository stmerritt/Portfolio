/// Header for SMERRITT
/// Clock Testbench Package

package vlab_clock_tb_pkg;
    // UVM library files
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "vlab_clock_tb_env.sv"
    `include "vlab_clock_tests.sv"
endpackage

